`timescale 1ns / 1ps

module vga_controller(
    input wire clk,
    input wire reset,
    output reg hsync,
    output reg vsync,
    output wire video_on,
    output wire [9:0] x,
    output wire [9:0] y
);

    parameter H_DISPLAY    = 640;
    parameter H_FRONT      = 16;
    parameter H_SYNC       = 96;
    parameter H_BACK       = 48;
    parameter H_TOTAL      = 800;

    parameter V_DISPLAY    = 480;
    parameter V_FRONT      = 10;
    parameter V_SYNC       = 2;
    parameter V_BACK       = 33;
    parameter V_TOTAL      = 525;

    reg [1:0] pixel_clk_count;
    reg pixel_clk;
    
    always @(posedge clk or posedge reset) begin
        if (reset) begin
            pixel_clk_count <= 0;
            pixel_clk <= 0;
        end else begin
            pixel_clk_count <= pixel_clk_count + 1;
            if (pixel_clk_count == 1) begin
                pixel_clk <= ~pixel_clk;
                pixel_clk_count <= 0;
            end
        end
    end

    reg [9:0] h_count;
    reg [9:0] v_count;

    always @(posedge pixel_clk or posedge reset) begin
        if (reset) begin
            h_count <= 0;
            v_count <= 0;
        end else begin
            if (h_count < H_TOTAL - 1) begin
                h_count <= h_count + 1;
            end else begin
                h_count <= 0;
                if (v_count < V_TOTAL - 1) begin
                    v_count <= v_count + 1;
                end else begin
                    v_count <= 0;
                end
            end
        end
    end

    always @(posedge pixel_clk or posedge reset) begin
        if (reset)
            hsync <= 1;
        else
            hsync <= (h_count >= (H_DISPLAY + H_FRONT)) && 
                     (h_count < (H_DISPLAY + H_FRONT + H_SYNC)) ? 0 : 1;
    end

    always @(posedge pixel_clk or posedge reset) begin
        if (reset)
            vsync <= 1;
        else
            vsync <= (v_count >= (V_DISPLAY + V_FRONT)) && 
                     (v_count < (V_DISPLAY + V_FRONT + V_SYNC)) ? 0 : 1;
    end

    assign video_on = (h_count < H_DISPLAY) && (v_count < V_DISPLAY);

    assign x = h_count;
    assign y = v_count;

endmodule